<?xml version="1.0" encoding="UTF-8"?>
<Batch version="2.0"><TaskList><Task type="ReplaceColorsTask" enabled="True"><FromType>0</FromType><FromColor>#717171</FromColor><FromTolerance>0</FromTolerance><FromColorStart>#808080</FromColorStart><FromColorEnd>#000000</FromColorEnd><FromAlphaStart>0</FromAlphaStart><FromAlphaEnd>255</FromAlphaEnd><ToType>0</ToType><ToColor>#91117E</ToColor><ToAlphaStart>0</ToAlphaStart><ToAlphaEnd>255</ToAlphaEnd></Task><Task type="ReplaceColorsTask" enabled="True"><FromType>0</FromType><FromColor>#404040</FromColor><FromTolerance>0</FromTolerance><FromColorStart>#808080</FromColorStart><FromColorEnd>#000000</FromColorEnd><FromAlphaStart>0</FromAlphaStart><FromAlphaEnd>255</FromAlphaEnd><ToType>0</ToType><ToColor>#2E1FCF</ToColor><ToAlphaStart>0</ToAlphaStart><ToAlphaEnd>255</ToAlphaEnd></Task><Task type="ReplaceColorsTask" enabled="True"><FromType>0</FromType><FromColor>#2D2D2D</FromColor><FromTolerance>0</FromTolerance><FromColorStart>#808080</FromColorStart><FromColorEnd>#000000</FromColorEnd><FromAlphaStart>0</FromAlphaStart><FromAlphaEnd>255</FromAlphaEnd><ToType>0</ToType><ToColor>#4A1212</ToColor><ToAlphaStart>0</ToAlphaStart><ToAlphaEnd>255</ToAlphaEnd></Task><Task type="ReplaceColorsTask" enabled="True"><FromType>0</FromType><FromColor>#D2D2D2</FromColor><FromTolerance>0</FromTolerance><FromColorStart>#808080</FromColorStart><FromColorEnd>#000000</FromColorEnd><FromAlphaStart>0</FromAlphaStart><FromAlphaEnd>255</FromAlphaEnd><ToType>0</ToType><ToColor>#E9D38C</ToColor><ToAlphaStart>0</ToAlphaStart><ToAlphaEnd>255</ToAlphaEnd></Task><Task type="ReplaceColorsTask" enabled="True"><FromType>0</FromType><FromColor>#969696</FromColor><FromTolerance>0</FromTolerance><FromColorStart>#808080</FromColorStart><FromColorEnd>#000000</FromColorEnd><FromAlphaStart>0</FromAlphaStart><FromAlphaEnd>255</FromAlphaEnd><ToType>0</ToType><ToColor>#751C0A</ToColor><ToAlphaStart>0</ToAlphaStart><ToAlphaEnd>255</ToAlphaEnd></Task><Task type="SaveAsTask" enabled="True"><FileName><![CDATA[Agent0003_<Original Name (Without Extension)>]]></FileName><PreserveStruct>False</PreserveStruct><CommonFolder><![CDATA[]]></CommonFolder><FileType></FileType><FilePath><![CDATA[D:\Workspace\IntelliJ\Serious Gaming\project\raw_assets\img\character\colored]]></FilePath><FileExists>0</FileExists><DefaultOptions>True</DefaultOptions><BMPCompression>0</BMPCompression><BMPVersion>1</BMPVersion><JPEGColorSpace>2</JPEGColorSpace><JPEGDCTMethod>0</JPEGDCTMethod><JPEGCromaSubsampling>1</JPEGCromaSubsampling><JPEGOptimalHuffman>False</JPEGOptimalHuffman><JPEGQuality>95</JPEGQuality><PNGCompression>5</PNGCompression><PNGFilter>1</PNGFilter><PNGInterlaced>False</PNGInterlaced><J2000ColorSpace>1</J2000ColorSpace><J2000Rate>0.500</J2000Rate><PCXCompression>1</PCXCompression><HDPLossless>False</HDPLossless><HDPImageQuality>0.900</HDPImageQuality><TGACompressed>False</TGACompressed><DDSMIPLevels>8</DDSMIPLevels><DDSMipMapFilter>4</DDSMipMapFilter><DDSFormat>71</DDSFormat><TIFFCompression>0</TIFFCompression><TIFFJPEGColorSpace>2</TIFFJPEGColorSpace><TIFFJPEGQuality>95</TIFFJPEGQuality><TIFFZIPCompression>1</TIFFZIPCompression><TIFFPlanarConf>1</TIFFPlanarConf><DICOMCompression>6</DICOMCompression><DICOMJPEG2000Rate>1</DICOMJPEG2000Rate><DICOMJPEGQuality>95</DICOMJPEGQuality></Task></TaskList></Batch>
